module vase

pub struct Updates {
	set string
	increment string
	append string
	prepend string
	delete string
}