module vase

pub struct Query {
	query string
	limit string
	last string
}